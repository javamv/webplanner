�� < d i v   c l a s s = " c o n t e n t L a y o u t 2 " > 
 < d i v   c l a s s = " c o l u m n L a y o u t   t w o - r i g h t - s i d e b a r "   d a t a - l a y o u t = " t w o - r i g h t - s i d e b a r " > 
 < d i v   c l a s s = " c e l l   n o r m a l "   d a t a - t y p e = " n o r m a l " > 
 < d i v   c l a s s = " i n n e r C e l l " > 
 	 < p > 
 	 	 < s p a n   s t y l e = " c o l o r :   r g b ( 1 0 2 , 1 0 2 , 1 0 2 ) ; " > 
 	 	 	 < s p a n   c l a s s = " c o n f l u e n c e - e m b e d d e d - f i l e - w r a p p e r   i m a g e - l e f t - w r a p p e r   c o n f l u e n c e - e m b e d d e d - m a n u a l - s i z e " > 
 	 	 	 	 < i m g   c l a s s = " c o n f l u e n c e - e m b e d d e d - i m a g e   c o n f l u e n c e - e x t e r n a l - r e s o u r c e   i m a g e - l e f t "   h e i g h t = " 2 5 0 "   s r c = " $ { i m a g e } "   d a t a - i m a g e - s r c = " $ { i m a g e } " / > 
 	 	 	 < / s p a n > 
 	 	 	 $ { d e s c r i p t i o n } 
 	 	 < / s p a n > 
 	 < / p > 
 	 < p > 
 	 	 < s p a n   c l a s s = " d e t a i l s "   s t y l e = " c o l o r :   r g b ( 1 0 2 , 1 0 2 , 1 0 2 ) ; " > & n b s p ; < / s p a n > 
 	 < / p > 
 	 < p > 
 	 	 < s t r o n g > < e m > T i m e < / e m > < / s t r o n g > 
 	 < / p > 
 	 < p > 
 	 	 < s p a n   c l a s s = " d e t a i l s "   s t y l e = " c o l o r :   r g b ( 1 0 2 , 1 0 2 , 1 0 2 ) ; " > $ { t i m e } < / s p a n > 
 	 < / p > 
 	 < p > 
 	 	 < s p a n   c l a s s = " d e t a i l s "   s t y l e = " c o l o r :   r g b ( 1 0 2 , 1 0 2 , 1 0 2 ) ; " > & n b s p ; < / s p a n > 
 	 < / p > 
 	 < p > 
 	 	 < s t r o n g > R e g i s t r a t i o n   < s p a n   c l a s s = " n o l i n k " > & n b s p ; < / s p a n > 
 	 	 < a   c l a s s = " e x t e r n a l - l i n k "   h r e f = " $ { g o t o L i n k } "   r e l = " n o f o l l o w " > 
 	 	 	 < s p a n   c l a s s = " n o l i n k " > R e g i s t r a t i o n   L i n k < / s p a n > 
 	 	 < / a > 
 	 	 < / s t r o n g > 
 	 < / p > 
 	 	 
 	 < p > < s p a n   c l a s s = " d e t a i l s "   s t y l e = " c o l o r :   r g b ( 1 0 2 , 1 0 2 , 1 0 2 ) ; " > < b r / > < / s p a n > < / p > 
 < / d i v > 
 < / d i v > 
 < d i v   c l a s s = " c e l l   a s i d e "   d a t a - t y p e = " a s i d e " > 
 < d i v   c l a s s = " i n n e r C e l l " > 
 < p > & n b s p ; < / p > < / d i v > 
 < / d i v > 
 < / d i v > 
 < / d i v >