�� < p > < s p a n   s t y l e = " c o l o r :   r g b ( 1 0 2 , 1 0 2 , 1 0 2 ) ; " > < s p a n   c l a s s = " c o n f l u e n c e - e m b e d d e d - f i l e - w r a p p e r   c o n f l u e n c e - e m b e d d e d - m a n u a l - s i z e " > < i m g   c l a s s = " c o n f l u e n c e - e m b e d d e d - i m a g e   c o n f l u e n c e - e x t e r n a l - r e s o u r c e "   h e i g h t = " 2 5 0 "   s r c = " $ { i m a g e } "   d a t a - i m a g e - s r c = " $ { i m a g e } " / > < / s p a n >   T h i s   w e b i n a r   a b o u t   n e w   a g i l e   m e t h o d s   < / s p a n > < / p >